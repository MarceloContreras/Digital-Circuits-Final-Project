library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Wallace8signed is
    Port ( a,b : in STD_LOGIC_VECTOR (7 downto 0);
           prod : out STD_LOGIC_VECTOR (15 downto 0));
end Wallace8signed;

architecture Behavioral of Wallace8signed is

begin


end Behavioral;
